library verilog;
use verilog.vl_types.all;
entity DX_reg_sv_unit is
end DX_reg_sv_unit;
