library verilog;
use verilog.vl_types.all;
entity MW_reg_sv_unit is
end MW_reg_sv_unit;
