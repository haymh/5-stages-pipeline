library verilog;
use verilog.vl_types.all;
entity FD_reg_sv_unit is
end FD_reg_sv_unit;
