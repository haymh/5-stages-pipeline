library verilog;
use verilog.vl_types.all;
entity XM_reg_sv_unit is
end XM_reg_sv_unit;
